module cache_ctrl();


endmodule